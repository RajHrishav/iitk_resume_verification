module prac_tb();
	
	reg [255:0] a, b;
	wire [511:0] prod;
	
	ks256 p(.a(a),.b(b),.prod(prod));
	
	initial 
		begin
			$monitor($time,"A = %b, B = %b, Y = %b",a,b,prod);
			// #5 a = 3'b111;b = 3'b111;
			//#5 a = 8'b00000111;b = 8'b00000001;
			//#5 a = 16'b0000000000001111;b = 16'b0000000000000010;
			//#5 a = 32'b0000000000000000000000000001111;b = 32'b0000000000000000000000000000010;
			//#5 a = 64'b00000000000000000000000000000000000000000000000000000000001111;b = 64'b00000000000000000000000000000000000000000000000000000000000010;
			#5 a = 256'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111;b = 256'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;
			#5 $finish;
		end
endmodule


